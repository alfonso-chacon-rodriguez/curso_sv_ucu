`ifndef DEFS_DONE
  `define DEFS_DONE //set the definitions done flag

  package definitions_pkg;

  parameter VERSION = "Curso-Uruguay-1.0";



endpackage

`endif

